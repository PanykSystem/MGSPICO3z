`ifndef DEFINES_SVH
`define DEFINES_SVH

`default_nettype none

`define	HIGH	1'b1
`define	LOW		1'b0

typedef	logic [21:0] psram_addr_t;

`default_nettype wire
`endif // DEFINES_SVH
