//`define IKASCC_SIMULATION
//`define IKASCC_ASYNC_VENDOR_ALTERA
//`define IKASCC_ASYNC_VENDOR_XILINX
//`define IKASCC_ASYNC_VENDOR_LATTICE
`define IKASCC_ASYNC_VENDOR_GOWIN
